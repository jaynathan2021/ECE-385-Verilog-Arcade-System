module score_text_rom
(
	input [7:0] address,
	output [7:0] data

);

	parameter[0:95][7:0] ROM = {

         // code x53
                8'b00000000, // 0  
                8'b00000000, // 1
                8'b11111110, // 2 *******
                8'b11111110, // 3  **  **
                8'b11000000, // 4  **   *
                8'b11000000, // 5  ** *
                8'b11111110, // 6  ****
                8'b11111110, // 7  ** *
                8'b00100100, // 8  **
                8'b00000110, // 9  **   *
                8'b11111110, // a  **  **
                8'b11111110, // b *******
                8'b00000000, // c
                8'b00000000, // d
                8'b00000000, // e
                8'b00000000, // f 

         // code x43
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111110, // 2   ****
        8'b11111110, // 3  **  **
        8'b11000010, // 4 **    *
        8'b11000000, // 5 **
        8'b11000000, // 6 **
        8'b11000000, // 7 **
        8'b11000000, // 8 **
        8'b11000010, // 9 **    *
        8'b11111110, // a  **  **
        8'b01111110, // b   ****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

         // code x4f
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111110, // 2  *****
        8'b11000110, // 3 **   **
        8'b11000110, // 4 **   **
        8'b11000110, // 5 **   **
        8'b11000110, // 6 **   **
        8'b11000110, // 7 **   **
        8'b11000110, // 8 **   **
        8'b11000110, // 9 **   **
        8'b11000110, // a **   **
        8'b11111110, // b  *****
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

         // code x52
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111110, // 2 ******
        8'b01111111, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01111111, // 6 *******
        8'b01111111, // 7 *******
        8'b01111100, // 8 **   **
        8'b01101110, // 9 **   **
        8'b01100111, // a **   **
        8'b01100111, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

         // code x45
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111111, // 2 *******
        8'b01111111, // 3 *******
        8'b01100000, // 4 **
        8'b01100000, // 5 **
        8'b01111111, // 6 *******
        8'b01111111, // 7 *******
        8'b01100000, // 8 **
        8'b01100000, // 9 **
        8'b01111111, // a *******
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
		  
         // code x3a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
	
	
	};
	
	assign data = ROM[address];

endmodule 



module score_text_map
(
	input logic [5:0] X,
	input logic [3:0] Y,
	output logic pixel
);

	logic [7:0] rom_address;
	logic [7:0] text_slice;
	
	assign pixel = text_slice[3'b111 - X[2:0]];

	score_text_rom text_rom(.address(rom_address), .data(text_slice));


	always_comb begin
	
		//S
		if(X >= 6'd0 && X < 6'd8) begin
			rom_address = 8'd0 + Y;
		end
		
		//C
		else if(X >= 6'd8 && X < 6'd16) begin
			rom_address = 8'd16 + Y;
		end
		
		//O
		else if(X >= 6'd16 && X < 6'd24) begin
			rom_address = 8'd32 + Y;
		end
		
		//R
		else if(X >= 6'd24 && X < 6'd32) begin
			rom_address = 8'd48 + Y;
		end
		
		//E
		else if(X >= 6'd32 && X < 6'd40) begin
			rom_address = 8'd64 + Y;
		end
		
		//:
		else begin
			rom_address = 8'd80 + Y;
		end
	
	end
	
endmodule 