module lives_text_rom
(
	input [7:0] address,
	output [7:0] data

);

	parameter[0:111][7:0] ROM = {
         // code x4c
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100011, // 2 **   **
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01111111, // 6 *******
        8'b01111111, // 7 *******
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b01100011, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

         // code x49
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01111111, // 2 *******
        8'b01111111, // 3 *******
        8'b01100000, // 4 **
        8'b01100000, // 5 **
        8'b01111111, // 6 *******
        8'b01111111, // 7 *******
        8'b01100000, // 8 **
        8'b01100000, // 9 **
        8'b01111111, // a *******
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
		  
         // code x56
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00111100, // 2   ****
        8'b01111110, // 3  ******
        8'b01100110, // 4  **  **
        8'b01100110, // 5  **  **
        8'b01111110, // 6  ******
        8'b01111110, // 7  ******
        8'b01100110, // 8  **  **
        8'b01100110, // 9  **  **
        8'b01100110, // a  **  **
        8'b01100110, // b  **  **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

         // code x45
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100000, // 2 **
        8'b01100000, // 3 **
        8'b01100000, // 4 **
        8'b01100000, // 5 **
        8'b01100000, // 6 **
        8'b01100000, // 7 **
        8'b01100000, // 8 **
        8'b01100000, // 9 **
        8'b01111111, // a *******
        8'b01111111, // b *******
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
		  
         // code x53
        8'b00000000, // 0
        8'b00000000, // 1
        8'b11111111, // 2 ********
        8'b11111111, // 3 ********
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00011000, // 6    **
        8'b00011000, // 7    **
        8'b00011000, // 8    **
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00011000, // b    **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f
		  
         // code x3a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b01100011, // 2 **   **
        8'b01100011, // 3 **   **
        8'b01100011, // 4 **   **
        8'b01100011, // 5 **   **
        8'b01111111, // 6 *******
        8'b01111111, // 7 *******
        8'b01100011, // 8 **   **
        8'b01100011, // 9 **   **
        8'b01100011, // a **   **
        8'b01100011, // b **   **
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f

	 // code x3a
        8'b00000000, // 0
        8'b00000000, // 1
        8'b00000000, // 2
        8'b00000000, // 3
        8'b00011000, // 4    **
        8'b00011000, // 5    **
        8'b00000000, // 6
        8'b00000000, // 7
        8'b00000000, // 8
        8'b00011000, // 9    **
        8'b00011000, // a    **
        8'b00000000, // b
        8'b00000000, // c
        8'b00000000, // d
        8'b00000000, // e
        8'b00000000, // f


	};
	
	assign data = ROM[address];

endmodule 

module lives_text_map
(
	input logic [5:0] X,
	input logic [3:0] Y,
	output logic pixel
);

	logic [7:0] rom_address;
	logic [7:0] text_slice;
	
	assign pixel = text_slice[3'b111 - X[2:0]];

	lives_text_rom text_rom(.address(rom_address), .data(text_slice));
	
	always_comb 
        begin
		
		//H
		if(X >= 6'd0 && X < 6'd8) begin
			rom_address = 8'd0 + Y;
		end
		
		//E
		else if(X >= 6'd8 && X < 6'd16) begin
			rom_address = 8'd16 + Y;
		end
		
		//A
		else if(X >= 6'd16 && X < 6'd24) begin
			rom_address = 8'd32 + Y;
		end
		
		//L
		else if(X >= 6'd24 && X < 6'd32) begin
			rom_address = 8'd48 + Y;
		end
		
		//T
		else if(X >= 6'd32 && X < 6'd40) begin
			rom_address = 8'd64 + Y;
		end
		//H
                else if(X >= 6'd40 && X < 6'd48) begin
			rom_address = 8'd80 + Y;
		end

		//:
		else begin
			rom_address = 8'd96 + Y;
		end
		
	end

endmodule 