module sprite_map(
						);
						
endmodule